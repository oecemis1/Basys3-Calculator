`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 13.08.2022 23:16:31
// Design Name: 
// Module Name: SevenSegmentDisplayer_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SevenSegmentDisplayer_tb(input clock_100Mhz);

    reg reset_tb;
    reg [6:0]whole_number_tb;
    reg [6:0]fraction_number;
    reg sign;
    



endmodule
